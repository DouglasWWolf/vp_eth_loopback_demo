//////////////////////////////////////
// ACE GENERATED VERILOG INCLUDE FILE
// Generated on: 2023.05.10 at 14:47:42 PDT
// By: ACE 9.0.1
// From project: vp_project
//////////////////////////////////////
// User Design Port Binding Include File
//////////////////////////////////////

//////////////////////////////////////
// User Design Ports
//////////////////////////////////////
    // Ports for ethernet_0
    // Clocks and Resets
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_m0_ff_clk_divby2, i_user_02_09_mt_00[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_m1_ff_clk_divby2, i_user_02_09_mt_00[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_ref_clk_divby2, i_user_02_09_mt_00[2])
    // Free Running Counter
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[0], o_user_02_09_lut_06[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[1], o_user_02_09_bram_01[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[2], o_user_02_09_bram_01[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[3], o_user_02_09_bram_01[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[4], o_user_02_09_bram_01[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[5], o_user_02_09_bram_01[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[6], o_user_02_09_bram_01[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[7], o_user_02_09_bram_01[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[8], o_user_02_09_bram_01[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[9], o_user_02_09_bram_01[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[10], o_user_02_09_bram_01[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[11], o_user_02_09_bram_01[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[12], o_user_02_09_bram_01[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[13], o_user_02_09_bram_01[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[14], o_user_02_09_bram_01[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[15], o_user_02_09_bram_01[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[16], o_user_02_09_bram_01[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[17], o_user_02_09_bram_01[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[18], o_user_02_09_bram_01[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[19], o_user_02_09_bram_01[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[20], o_user_02_09_bram_01[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[21], o_user_02_09_bram_01[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[22], o_user_02_09_bram_01[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[23], o_user_02_09_mlp_01[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[24], o_user_02_09_mlp_01[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[25], o_user_02_09_mlp_01[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[26], o_user_02_09_mlp_01[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[27], o_user_02_09_mlp_01[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[28], o_user_02_09_mlp_01[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[29], o_user_02_09_mlp_01[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[30], o_user_02_09_mlp_01[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[31], o_user_02_09_mlp_01[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[32], o_user_02_09_mlp_01[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[33], o_user_02_09_mlp_01[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[34], o_user_02_09_mlp_01[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[35], o_user_02_09_mlp_01[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[36], o_user_02_09_mlp_01[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[37], o_user_02_09_mlp_01[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[38], o_user_02_09_mlp_01[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[39], o_user_02_09_mlp_01[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[40], o_user_02_09_mlp_01[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[41], o_user_02_09_mlp_01[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[42], o_user_02_09_mlp_01[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[43], o_user_02_09_mlp_01[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[44], o_user_02_09_mlp_01[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[45], o_user_02_09_mlp_01[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[46], o_user_02_09_lut_07[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[47], o_user_02_09_lut_07[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[48], o_user_02_09_lut_07[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[49], o_user_02_09_lut_07[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[50], o_user_02_09_lut_07[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[51], o_user_02_09_lut_07[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[52], o_user_02_09_lut_07[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[53], o_user_02_09_lut_07[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[54], o_user_02_09_lut_07[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[55], o_user_02_09_lut_07[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[56], o_user_02_09_lut_07[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[57], o_user_02_09_lut_07[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[58], o_user_02_09_lut_07[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[59], o_user_02_09_lut_07[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[60], o_user_02_09_lut_07[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[61], o_user_02_09_lut_07[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[62], o_user_02_09_lut_07[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_free_running_counter[63], o_user_02_09_lut_07[22])
    // Quad MAC 0 Flow Control
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_enable[0], i_user_02_09_lut_18[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_enable[1], i_user_02_09_lut_18[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_enable[2], i_user_02_09_lut_18[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_enable[3], i_user_02_09_lut_18[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_en[0], i_user_02_09_lut_17[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_en[1], i_user_02_09_lut_17[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_en[2], i_user_02_09_lut_17[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_en[3], i_user_02_09_lut_17[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[0], i_user_02_09_mlp_03[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[1], i_user_02_09_lut_16[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[2], i_user_02_09_lut_16[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[3], i_user_02_09_lut_16[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[4], i_user_02_09_lut_16[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[5], i_user_02_09_lut_16[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[6], i_user_02_09_lut_16[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[7], i_user_02_09_lut_16[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[8], i_user_02_09_lut_16[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[9], i_user_02_09_lut_16[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[10], i_user_02_09_lut_16[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[11], i_user_02_09_lut_16[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[12], i_user_02_09_lut_16[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[13], i_user_02_09_lut_16[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[14], i_user_02_09_lut_16[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[15], i_user_02_09_lut_16[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[16], i_user_02_09_lut_16[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[17], i_user_02_09_lut_16[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[18], i_user_02_09_lut_16[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[19], i_user_02_09_lut_16[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[20], i_user_02_09_lut_16[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[21], i_user_02_09_lut_17[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[22], i_user_02_09_lut_17[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[23], i_user_02_09_lut_17[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[24], i_user_02_09_lut_17[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[25], i_user_02_09_lut_17[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[26], i_user_02_09_lut_17[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[27], i_user_02_09_lut_17[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[28], i_user_02_09_lut_17[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[29], i_user_02_09_lut_17[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[30], i_user_02_09_lut_17[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_pause_on[31], i_user_02_09_lut_17[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[0], o_user_02_09_lut_16[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[1], o_user_02_09_lut_16[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[2], o_user_02_09_lut_16[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[3], o_user_02_09_lut_16[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[4], o_user_02_09_lut_16[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[5], o_user_02_09_lut_16[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[6], o_user_02_09_lut_16[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[7], o_user_02_09_lut_16[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[8], o_user_02_09_lut_16[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[9], o_user_02_09_lut_16[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[10], o_user_02_09_lut_16[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[11], o_user_02_09_lut_16[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[12], o_user_02_09_lut_16[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[13], o_user_02_09_lut_16[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[14], o_user_02_09_lut_16[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[15], o_user_02_09_lut_16[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[16], o_user_02_09_lut_16[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[17], o_user_02_09_lut_17[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[18], o_user_02_09_lut_17[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[19], o_user_02_09_lut_17[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[20], o_user_02_09_lut_17[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[21], o_user_02_09_lut_17[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[22], o_user_02_09_lut_17[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[23], o_user_02_09_lut_17[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[24], o_user_02_09_lut_17[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[25], o_user_02_09_lut_17[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[26], o_user_02_09_lut_17[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[27], o_user_02_09_lut_17[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[28], o_user_02_09_lut_17[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[29], o_user_02_09_lut_17[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[30], o_user_02_09_lut_17[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_emac_xoff_gen[31], o_user_02_09_lut_17[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_lpi_txhold[0], o_user_02_09_lut_18[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_lpi_txhold[1], o_user_02_09_lut_18[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_lpi_txhold[2], o_user_02_09_lut_18[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_lpi_txhold[3], o_user_02_09_lut_18[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_mac_stop_tx[0], o_user_02_09_lut_17[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_mac_stop_tx[1], o_user_02_09_lut_17[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_mac_stop_tx[2], o_user_02_09_lut_17[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_mac_stop_tx[3], o_user_02_09_lut_17[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_hold_req[0], o_user_02_09_lut_18[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_hold_req[1], o_user_02_09_lut_18[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_hold_req[2], o_user_02_09_lut_18[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_hold_req[3], o_user_02_09_lut_18[9])
    // Quad MAC 0 Status
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_m0_ffe_tx_ovr[0], i_user_02_09_lut_18[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_m0_ffe_tx_ovr[1], i_user_02_09_lut_18[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_m0_ffe_tx_ovr[2], i_user_02_09_lut_18[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_m0_ffe_tx_ovr[3], i_user_02_09_lut_18[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_m0_ffp_tx_ovr[0], i_user_02_09_lut_18[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_m0_ffp_tx_ovr[1], i_user_02_09_lut_18[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_m0_ffp_tx_ovr[2], i_user_02_09_lut_18[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_m0_ffp_tx_ovr[3], i_user_02_09_lut_18[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_m0_mac_tx_underflow[0], i_user_02_09_lut_18[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_m0_mac_tx_underflow[1], i_user_02_09_lut_18[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_m0_mac_tx_underflow[2], i_user_02_09_lut_18[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_m0_mac_tx_underflow[3], i_user_02_09_lut_18[24])
    // Quad MAC 0 TSN
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[0], i_user_02_09_lut_05[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[1], i_user_02_09_lut_05[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[2], i_user_02_09_lut_05[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[3], i_user_02_09_lut_05[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[4], i_user_02_09_lut_05[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[5], i_user_02_09_lut_05[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[6], i_user_02_09_lut_05[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[7], i_user_02_09_lut_05[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[8], i_user_02_09_lut_05[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[9], i_user_02_09_lut_06[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[10], i_user_02_09_lut_06[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[11], i_user_02_09_lut_06[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[12], i_user_02_09_lut_06[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[13], i_user_02_09_lut_06[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[14], i_user_02_09_lut_06[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[15], i_user_02_09_lut_06[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[16], i_user_02_09_lut_06[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[17], i_user_02_09_lut_06[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[18], i_user_02_09_lut_06[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[19], i_user_02_09_lut_06[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[20], i_user_02_09_lut_06[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[21], i_user_02_09_lut_06[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[22], i_user_02_09_lut_06[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[23], i_user_02_09_lut_06[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[24], i_user_02_09_lut_06[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[25], i_user_02_09_lut_06[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[26], i_user_02_09_lut_06[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[27], i_user_02_09_lut_06[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[28], i_user_02_09_lut_06[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[29], i_user_02_09_lut_06[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[30], i_user_02_09_lut_06[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[31], i_user_02_09_lut_06[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[32], i_user_02_09_bram_01[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[33], i_user_02_09_bram_01[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[34], i_user_02_09_bram_01[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[35], i_user_02_09_bram_01[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[36], i_user_02_09_bram_01[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[37], i_user_02_09_bram_01[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[38], i_user_02_09_bram_01[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[39], i_user_02_09_bram_01[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[40], i_user_02_09_bram_01[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[41], i_user_02_09_bram_01[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[42], i_user_02_09_bram_01[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[43], i_user_02_09_bram_01[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[44], i_user_02_09_bram_01[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[45], i_user_02_09_bram_01[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[46], i_user_02_09_bram_01[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[47], i_user_02_09_bram_01[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[48], i_user_02_09_bram_01[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[49], i_user_02_09_bram_01[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[50], i_user_02_09_bram_01[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[51], i_user_02_09_bram_01[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[52], i_user_02_09_bram_01[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[53], i_user_02_09_bram_01[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[54], i_user_02_09_mlp_01[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[55], i_user_02_09_mlp_01[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[56], i_user_02_09_mlp_01[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[57], i_user_02_09_mlp_01[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[58], i_user_02_09_mlp_01[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[59], i_user_02_09_mlp_01[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[60], i_user_02_09_mlp_01[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[61], i_user_02_09_mlp_01[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[62], i_user_02_09_mlp_01[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[63], i_user_02_09_mlp_01[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[64], i_user_02_09_mlp_01[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[65], i_user_02_09_mlp_01[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[66], i_user_02_09_mlp_01[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[67], i_user_02_09_mlp_01[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[68], i_user_02_09_mlp_01[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[69], i_user_02_09_mlp_01[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[70], i_user_02_09_mlp_01[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[71], i_user_02_09_mlp_01[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[72], i_user_02_09_mlp_01[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[73], i_user_02_09_mlp_01[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[74], i_user_02_09_mlp_01[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[75], i_user_02_09_mlp_01[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[76], i_user_02_09_mlp_01[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[77], i_user_02_09_lut_07[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[78], i_user_02_09_lut_07[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[79], i_user_02_09_lut_07[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[80], i_user_02_09_lut_07[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[81], i_user_02_09_lut_07[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[82], i_user_02_09_lut_07[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[83], i_user_02_09_lut_07[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[84], i_user_02_09_lut_07[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[85], i_user_02_09_lut_07[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[86], i_user_02_09_lut_07[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[87], i_user_02_09_lut_07[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[88], i_user_02_09_lut_07[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[89], i_user_02_09_lut_07[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[90], i_user_02_09_lut_07[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[91], i_user_02_09_lut_07[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[92], i_user_02_09_lut_07[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[93], i_user_02_09_lut_07[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[94], i_user_02_09_lut_07[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[95], i_user_02_09_lut_07[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[96], i_user_02_09_lut_07[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[97], i_user_02_09_lut_07[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[98], i_user_02_09_lut_07[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[99], i_user_02_09_lut_08[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[100], i_user_02_09_lut_08[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[101], i_user_02_09_lut_08[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[102], i_user_02_09_lut_08[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[103], i_user_02_09_lut_08[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[104], i_user_02_09_lut_08[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[105], i_user_02_09_lut_08[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[106], i_user_02_09_lut_08[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[107], i_user_02_09_lut_08[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[108], i_user_02_09_lut_08[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[109], i_user_02_09_lut_08[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[110], i_user_02_09_lut_08[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[111], i_user_02_09_lut_08[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[112], i_user_02_09_lut_08[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[113], i_user_02_09_lut_08[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[114], i_user_02_09_lut_08[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[115], i_user_02_09_lut_08[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[116], i_user_02_09_lut_08[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[117], i_user_02_09_lut_08[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[118], i_user_02_09_lut_08[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[119], i_user_02_09_lut_08[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[120], i_user_02_09_lut_08[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[121], i_user_02_09_lut_08[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[122], i_user_02_09_lut_09[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[123], i_user_02_09_lut_09[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[124], i_user_02_09_lut_09[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[125], i_user_02_09_lut_09[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[126], i_user_02_09_lut_09[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[127], i_user_02_09_lut_09[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[128], i_user_02_09_lut_00[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[129], i_user_02_09_lut_01[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[130], i_user_02_09_lut_01[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[131], i_user_02_09_lut_01[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[132], i_user_02_09_lut_01[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[133], i_user_02_09_lut_01[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[134], i_user_02_09_lut_01[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[135], i_user_02_09_lut_01[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[136], i_user_02_09_lut_01[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[137], i_user_02_09_lut_01[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[138], i_user_02_09_lut_01[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[139], i_user_02_09_lut_01[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[140], i_user_02_09_lut_01[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[141], i_user_02_09_lut_01[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[142], i_user_02_09_lut_01[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[143], i_user_02_09_lut_01[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[144], i_user_02_09_lut_01[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[145], i_user_02_09_lut_01[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[146], i_user_02_09_lut_01[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[147], i_user_02_09_lut_01[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[148], i_user_02_09_lut_01[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[149], i_user_02_09_lut_01[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[150], i_user_02_09_lut_01[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[151], i_user_02_09_lut_01[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[152], i_user_02_09_lut_02[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[153], i_user_02_09_lut_02[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[154], i_user_02_09_lut_02[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[155], i_user_02_09_lut_02[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[156], i_user_02_09_lut_02[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[157], i_user_02_09_lut_02[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[158], i_user_02_09_lut_02[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[159], i_user_02_09_lut_02[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[160], i_user_02_09_lut_02[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[161], i_user_02_09_lut_02[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[162], i_user_02_09_lut_02[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[163], i_user_02_09_lut_02[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[164], i_user_02_09_lut_02[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[165], i_user_02_09_lut_02[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[166], i_user_02_09_lut_02[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[167], i_user_02_09_lut_02[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[168], i_user_02_09_lut_02[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[169], i_user_02_09_lut_02[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[170], i_user_02_09_lut_02[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[171], i_user_02_09_lut_02[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[172], i_user_02_09_lut_02[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[173], i_user_02_09_lut_02[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[174], i_user_02_09_bram_00[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[175], i_user_02_09_bram_00[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[176], i_user_02_09_bram_00[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[177], i_user_02_09_bram_00[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[178], i_user_02_09_bram_00[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[179], i_user_02_09_bram_00[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[180], i_user_02_09_bram_00[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[181], i_user_02_09_bram_00[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[182], i_user_02_09_bram_00[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[183], i_user_02_09_bram_00[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[184], i_user_02_09_bram_00[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[185], i_user_02_09_bram_00[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[186], i_user_02_09_bram_00[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[187], i_user_02_09_bram_00[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[188], i_user_02_09_bram_00[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[189], i_user_02_09_bram_00[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[190], i_user_02_09_bram_00[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[191], i_user_02_09_bram_00[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[192], i_user_02_09_bram_00[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[193], i_user_02_09_bram_00[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[194], i_user_02_09_bram_00[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[195], i_user_02_09_bram_00[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[196], i_user_02_09_bram_00[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[197], i_user_02_09_mlp_00[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[198], i_user_02_09_mlp_00[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[199], i_user_02_09_mlp_00[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[200], i_user_02_09_mlp_00[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[201], i_user_02_09_mlp_00[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[202], i_user_02_09_mlp_00[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[203], i_user_02_09_mlp_00[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[204], i_user_02_09_mlp_00[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[205], i_user_02_09_mlp_00[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[206], i_user_02_09_mlp_00[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[207], i_user_02_09_mlp_00[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[208], i_user_02_09_mlp_00[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[209], i_user_02_09_mlp_00[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[210], i_user_02_09_mlp_00[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[211], i_user_02_09_mlp_00[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[212], i_user_02_09_mlp_00[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[213], i_user_02_09_mlp_00[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[214], i_user_02_09_mlp_00[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[215], i_user_02_09_mlp_00[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[216], i_user_02_09_mlp_00[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[217], i_user_02_09_mlp_00[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[218], i_user_02_09_mlp_00[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[219], i_user_02_09_lut_03[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[220], i_user_02_09_lut_03[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[221], i_user_02_09_lut_03[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[222], i_user_02_09_lut_03[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[223], i_user_02_09_lut_03[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[224], i_user_02_09_lut_03[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[225], i_user_02_09_lut_03[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[226], i_user_02_09_lut_03[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[227], i_user_02_09_lut_03[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[228], i_user_02_09_lut_03[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[229], i_user_02_09_lut_03[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[230], i_user_02_09_lut_03[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[231], i_user_02_09_lut_03[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[232], i_user_02_09_lut_03[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[233], i_user_02_09_lut_03[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[234], i_user_02_09_lut_03[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[235], i_user_02_09_lut_03[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[236], i_user_02_09_lut_03[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[237], i_user_02_09_lut_03[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[238], i_user_02_09_lut_03[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[239], i_user_02_09_lut_03[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[240], i_user_02_09_lut_03[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[241], i_user_02_09_lut_04[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[242], i_user_02_09_lut_04[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[243], i_user_02_09_lut_04[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[244], i_user_02_09_lut_04[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[245], i_user_02_09_lut_04[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[246], i_user_02_09_lut_04[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[247], i_user_02_09_lut_04[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[248], i_user_02_09_lut_04[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[249], i_user_02_09_lut_04[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[250], i_user_02_09_lut_04[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[251], i_user_02_09_lut_04[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[252], i_user_02_09_lut_04[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[253], i_user_02_09_lut_04[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[254], i_user_02_09_lut_04[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts[255], i_user_02_09_lut_04[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[0], i_user_02_09_lut_12[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[1], i_user_02_09_lut_12[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[2], i_user_02_09_lut_12[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[3], i_user_02_09_lut_12[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[4], i_user_02_09_lut_12[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[5], i_user_02_09_lut_12[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[6], i_user_02_09_lut_12[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[7], i_user_02_09_lut_12[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[8], i_user_02_09_lut_12[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[9], i_user_02_09_lut_12[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[10], i_user_02_09_lut_12[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[11], i_user_02_09_lut_12[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[12], i_user_02_09_lut_12[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[13], i_user_02_09_lut_12[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[14], i_user_02_09_lut_12[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_id[15], i_user_02_09_lut_12[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_val[0], i_user_02_09_lut_12[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_val[1], i_user_02_09_lut_12[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_val[2], i_user_02_09_lut_12[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_tx_ts_val[3], i_user_02_09_lut_12[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[0], o_user_02_09_lut_10[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[1], o_user_02_09_lut_10[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[2], o_user_02_09_lut_10[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[3], o_user_02_09_lut_10[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[4], o_user_02_09_lut_10[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[5], o_user_02_09_lut_10[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[6], o_user_02_09_lut_10[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[7], o_user_02_09_lut_10[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[8], o_user_02_09_lut_10[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[9], o_user_02_09_lut_10[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[10], o_user_02_09_lut_10[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[11], o_user_02_09_lut_10[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[12], o_user_02_09_lut_10[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[13], o_user_02_09_bram_02[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[14], o_user_02_09_bram_02[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[15], o_user_02_09_bram_02[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[16], o_user_02_09_bram_02[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[17], o_user_02_09_bram_02[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[18], o_user_02_09_bram_02[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[19], o_user_02_09_bram_02[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[20], o_user_02_09_bram_02[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[21], o_user_02_09_bram_02[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[22], o_user_02_09_bram_02[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[23], o_user_02_09_bram_02[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[24], o_user_02_09_bram_02[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[25], o_user_02_09_bram_02[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[26], o_user_02_09_bram_02[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[27], o_user_02_09_bram_02[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[28], o_user_02_09_bram_02[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[29], o_user_02_09_bram_02[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[30], o_user_02_09_bram_02[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[31], o_user_02_09_bram_02[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[32], o_user_02_09_bram_02[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[33], o_user_02_09_bram_02[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[34], o_user_02_09_bram_02[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[35], o_user_02_09_mlp_02[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[36], o_user_02_09_mlp_02[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[37], o_user_02_09_mlp_02[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[38], o_user_02_09_mlp_02[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[39], o_user_02_09_mlp_02[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[40], o_user_02_09_mlp_02[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[41], o_user_02_09_mlp_02[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[42], o_user_02_09_mlp_02[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[43], o_user_02_09_mlp_02[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[44], o_user_02_09_mlp_02[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[45], o_user_02_09_mlp_02[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[46], o_user_02_09_mlp_02[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[47], o_user_02_09_mlp_02[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[48], o_user_02_09_mlp_02[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[49], o_user_02_09_mlp_02[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[50], o_user_02_09_mlp_02[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[51], o_user_02_09_mlp_02[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[52], o_user_02_09_mlp_02[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[53], o_user_02_09_mlp_02[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[54], o_user_02_09_mlp_02[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[55], o_user_02_09_mlp_02[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[56], o_user_02_09_mlp_02[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[57], o_user_02_09_lut_11[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[58], o_user_02_09_lut_11[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[59], o_user_02_09_lut_11[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[60], o_user_02_09_lut_11[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[61], o_user_02_09_lut_11[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[62], o_user_02_09_lut_11[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[63], o_user_02_09_lut_11[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[64], o_user_02_09_lut_11[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[65], o_user_02_09_lut_11[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[66], o_user_02_09_lut_11[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[67], o_user_02_09_lut_11[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[68], o_user_02_09_lut_11[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[69], o_user_02_09_lut_11[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[70], o_user_02_09_lut_11[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[71], o_user_02_09_lut_11[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[72], o_user_02_09_lut_11[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[73], o_user_02_09_lut_11[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[74], o_user_02_09_lut_11[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[75], o_user_02_09_lut_11[22])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[76], o_user_02_09_lut_11[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[77], o_user_02_09_lut_11[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[78], o_user_02_09_lut_11[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[79], o_user_02_09_lut_11[27])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[80], o_user_02_09_lut_12[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[81], o_user_02_09_lut_12[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[82], o_user_02_09_lut_12[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[83], o_user_02_09_lut_12[4])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[84], o_user_02_09_lut_12[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[85], o_user_02_09_lut_12[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[86], o_user_02_09_lut_12[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[87], o_user_02_09_lut_12[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[88], o_user_02_09_lut_12[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[89], o_user_02_09_lut_12[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[90], o_user_02_09_lut_12[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[91], o_user_02_09_lut_12[14])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[92], o_user_02_09_lut_12[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[93], o_user_02_09_lut_12[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[94], o_user_02_09_lut_12[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[95], o_user_02_09_lut_12[19])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[96], o_user_02_09_lut_12[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[97], o_user_02_09_lut_12[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[98], o_user_02_09_lut_12[23])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[99], o_user_02_09_lut_12[24])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[100], o_user_02_09_lut_12[25])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[101], o_user_02_09_lut_12[26])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[102], o_user_02_09_lut_13[0])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[103], o_user_02_09_lut_13[1])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[104], o_user_02_09_lut_13[2])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[105], o_user_02_09_lut_13[3])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[106], o_user_02_09_lut_13[5])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[107], o_user_02_09_lut_13[6])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[108], o_user_02_09_lut_13[7])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[109], o_user_02_09_lut_13[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[110], o_user_02_09_lut_13[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[111], o_user_02_09_lut_13[11])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[112], o_user_02_09_lut_13[12])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[113], o_user_02_09_lut_13[13])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[114], o_user_02_09_lut_13[15])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[115], o_user_02_09_lut_13[16])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[116], o_user_02_09_lut_13[17])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[117], o_user_02_09_lut_13[18])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[118], o_user_02_09_lut_13[20])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay[119], o_user_02_09_lut_13[21])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay_val[0], o_user_02_09_lut_10[8])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay_val[1], o_user_02_09_lut_10[9])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay_val[2], o_user_02_09_lut_10[10])
`ACX_BIND_USER_DESIGN_PORT(ethernet_0_quad0_peer_delay_val[3], o_user_02_09_lut_10[11])
    // Ports for noc
    // Ports for pll_ddr
`ifdef ACX_CLK_SW_FULL
`ACX_BIND_USER_DESIGN_PORT(pll_ddr_lock, i_user_00_01_lut_17[0])
`endif
    // Ports for pll_eth_sys_ne_0
`ifdef ACX_CLK_NE_FULL
`ACX_BIND_USER_DESIGN_PORT(pll_eth_sys_ne_0_lock, i_user_12_08_lut_17[0])
`endif
    // Ports for pll_gddr_SE
`ifdef ACX_CLK_SE_FULL
`ACX_BIND_USER_DESIGN_PORT(pll_gddr_SE_lock, i_user_12_01_lut_17[0])
`endif
    // Ports for pll_gddr_SW
`ifdef ACX_CLK_SW_FULL
`ACX_BIND_USER_DESIGN_PORT(pll_gddr_SW_lock, i_user_00_01_lut_17[1])
`endif
    // Ports for pll_noc_ne_1
`ifdef ACX_CLK_NE_FULL
`ACX_BIND_USER_DESIGN_PORT(i_clk, i_user_06_09_trunk_00[21])
`ACX_BIND_USER_DESIGN_PORT(i_eth_ts_clk, i_user_06_09_trunk_00[20])
`ACX_BIND_USER_DESIGN_PORT(i_reg_clk, i_user_06_09_trunk_00[19])
`ACX_BIND_USER_DESIGN_PORT(pll_noc_ne_1_lock, i_user_12_08_lut_17[1])
`endif
    // Ports for pll_pcie
`ifdef ACX_CLK_NE_FULL
`ACX_BIND_USER_DESIGN_PORT(pll_pcie_lock, i_user_12_08_lut_17[2])
`endif
    // Ports for vp_clkio_ne
`ACX_BIND_USER_DESIGN_PORT(fpga_rst_l, i_user_06_09_trunk_00[127])
    // Ports for vp_clkio_nw
    // Ports for vp_clkio_se
    // Ports for vp_clkio_sw
    // Ports for vp_gpio_n_b0
`ifdef ACX_GPIO_N_FULL
    // Core Data
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_in[0], i_user_11_09_lut_13[15])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_in[1], i_user_11_09_lut_13[23])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_in[2], i_user_11_09_lut_14[3])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_in[3], i_user_11_09_lut_14[11])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_in[4], i_user_11_09_lut_14[19])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_in[5], i_user_11_09_lut_14[27])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_in[6], i_user_11_09_lut_15[7])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_in[7], i_user_11_09_lut_15[15])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_oe[0], o_user_11_09_lut_12[16])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_oe[1], o_user_11_09_lut_12[17])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_oe[2], o_user_11_09_lut_12[18])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_oe[3], o_user_11_09_lut_12[19])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_oe[4], o_user_11_09_lut_12[20])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_oe[5], o_user_11_09_lut_12[21])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_oe[6], o_user_11_09_lut_12[22])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_oe[7], o_user_11_09_lut_12[23])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_out[0], o_user_11_09_lut_13[12])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_out[1], o_user_11_09_lut_13[20])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_out[2], o_user_11_09_lut_14[0])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_out[3], o_user_11_09_lut_14[8])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_out[4], o_user_11_09_lut_14[16])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_out[5], o_user_11_09_lut_14[24])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_out[6], o_user_11_09_lut_15[4])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_fpga_out[7], o_user_11_09_lut_15[12])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_oe_l, o_user_11_09_lut_12[24])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_oe_l_oe, o_user_11_09_lut_12[14])
`ACX_BIND_USER_DESIGN_PORT(led_oe_l, o_user_11_09_lut_13[4])
`ACX_BIND_USER_DESIGN_PORT(led_oe_l_oe, o_user_11_09_lut_12[15])
`endif
    // Ports for vp_gpio_n_b1
`ifdef ACX_GPIO_N_FULL
    // Core Data
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir[0], o_user_11_09_lut_10[6])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir[1], o_user_11_09_lut_10[14])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir[2], o_user_11_09_lut_10[22])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir[3], o_user_11_09_lut_11[2])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir[4], o_user_11_09_lut_11[10])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir[5], o_user_11_09_lut_11[18])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir[6], o_user_11_09_lut_11[26])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir[7], o_user_11_09_lut_12[6])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir_oe[0], o_user_11_09_lut_09[10])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir_oe[1], o_user_11_09_lut_09[11])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir_oe[2], o_user_11_09_lut_09[12])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir_oe[3], o_user_11_09_lut_09[13])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir_oe[4], o_user_11_09_lut_09[14])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir_oe[5], o_user_11_09_lut_09[15])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir_oe[6], o_user_11_09_lut_09[16])
`ACX_BIND_USER_DESIGN_PORT(ext_gpio_dir_oe[7], o_user_11_09_lut_09[17])
`ACX_BIND_USER_DESIGN_PORT(led_l[4], o_user_11_09_lut_09[18])
`ACX_BIND_USER_DESIGN_PORT(led_l[5], o_user_11_09_lut_09[26])
`ACX_BIND_USER_DESIGN_PORT(led_l_oe[4], o_user_11_09_lut_09[8])
`ACX_BIND_USER_DESIGN_PORT(led_l_oe[5], o_user_11_09_lut_09[9])
`endif
    // Ports for vp_gpio_n_b2
`ifdef ACX_GPIO_N_FULL
    // Core Data
`ACX_BIND_USER_DESIGN_PORT(led_l[0], o_user_11_09_lut_07[0])
`ACX_BIND_USER_DESIGN_PORT(led_l[1], o_user_11_09_lut_07[8])
`ACX_BIND_USER_DESIGN_PORT(led_l[2], o_user_11_09_lut_07[16])
`ACX_BIND_USER_DESIGN_PORT(led_l[3], o_user_11_09_lut_07[24])
`ACX_BIND_USER_DESIGN_PORT(led_l[6], o_user_11_09_lut_08[4])
`ACX_BIND_USER_DESIGN_PORT(led_l[7], o_user_11_09_lut_08[12])
`ACX_BIND_USER_DESIGN_PORT(led_l_oe[0], o_user_11_09_lut_06[4])
`ACX_BIND_USER_DESIGN_PORT(led_l_oe[1], o_user_11_09_lut_06[5])
`ACX_BIND_USER_DESIGN_PORT(led_l_oe[2], o_user_11_09_lut_06[6])
`ACX_BIND_USER_DESIGN_PORT(led_l_oe[3], o_user_11_09_lut_06[7])
`ACX_BIND_USER_DESIGN_PORT(led_l_oe[6], o_user_11_09_lut_06[8])
`ACX_BIND_USER_DESIGN_PORT(led_l_oe[7], o_user_11_09_lut_06[9])
`endif
    // Ports for vp_gpio_s_b0
`ifdef ACX_GPIO_S_FULL
    // Core Data
`ACX_BIND_USER_DESIGN_PORT(fpga_avr_rxd, i_user_10_00_lut_07[7])
`ACX_BIND_USER_DESIGN_PORT(fpga_ftdi_rxd, i_user_10_00_lut_07[23])
`ACX_BIND_USER_DESIGN_PORT(fpga_i2c_mux_gnt, i_user_10_00_lut_06[11])
`ACX_BIND_USER_DESIGN_PORT(irq_to_fpga, i_user_10_00_lut_08[3])
`ACX_BIND_USER_DESIGN_PORT(qsfp_int_fpga_l, i_user_10_00_lut_06[3])
`ACX_BIND_USER_DESIGN_PORT(fpga_avr_txd, o_user_10_00_lut_07[26])
`ACX_BIND_USER_DESIGN_PORT(fpga_avr_txd_oe, o_user_10_00_lut_06[16])
`ACX_BIND_USER_DESIGN_PORT(fpga_ftdi_txd, o_user_10_00_lut_08[14])
`ACX_BIND_USER_DESIGN_PORT(fpga_ftdi_txd_oe, o_user_10_00_lut_06[18])
`ACX_BIND_USER_DESIGN_PORT(fpga_i2c_req_l, o_user_10_00_lut_07[18])
`ACX_BIND_USER_DESIGN_PORT(fpga_i2c_req_l_oe, o_user_10_00_lut_06[15])
`ACX_BIND_USER_DESIGN_PORT(irq_to_avr, o_user_10_00_lut_09[10])
`ACX_BIND_USER_DESIGN_PORT(irq_to_avr_oe, o_user_10_00_lut_06[21])
`ACX_BIND_USER_DESIGN_PORT(test[1], o_user_10_00_lut_06[22])
`ACX_BIND_USER_DESIGN_PORT(test_oe[1], o_user_10_00_lut_06[12])
`endif
    // Ports for vp_gpio_s_b1
`ifdef ACX_GPIO_S_FULL
    // Core Clock
`ACX_BIND_USER_DESIGN_PORT(mcio_vio_45_10_clk, i_user_10_00_mt_00[1])
    // Core Data
`ACX_BIND_USER_DESIGN_PORT(mcio_vio_in[0], i_user_10_00_lut_03[14])
`ACX_BIND_USER_DESIGN_PORT(mcio_vio_in[1], i_user_10_00_lut_03[22])
`ACX_BIND_USER_DESIGN_PORT(mcio_vio_in[2], i_user_10_00_lut_04[2])
`ACX_BIND_USER_DESIGN_PORT(mcio_vio_in[3], i_user_10_00_lut_04[10])
`ACX_BIND_USER_DESIGN_PORT(mcio_dir[0], o_user_10_00_lut_05[8])
`ACX_BIND_USER_DESIGN_PORT(mcio_dir[1], o_user_10_00_lut_05[16])
`ACX_BIND_USER_DESIGN_PORT(mcio_dir[2], o_user_10_00_lut_05[24])
`ACX_BIND_USER_DESIGN_PORT(mcio_dir[3], o_user_10_00_lut_06[4])
`ACX_BIND_USER_DESIGN_PORT(mcio_dir_45, o_user_10_00_lut_03[16])
`ACX_BIND_USER_DESIGN_PORT(mcio_dir_45_oe, o_user_10_00_lut_03[6])
`ACX_BIND_USER_DESIGN_PORT(mcio_dir_oe[0], o_user_10_00_lut_03[12])
`ACX_BIND_USER_DESIGN_PORT(mcio_dir_oe[1], o_user_10_00_lut_03[13])
`ACX_BIND_USER_DESIGN_PORT(mcio_dir_oe[2], o_user_10_00_lut_03[14])
`ACX_BIND_USER_DESIGN_PORT(mcio_dir_oe[3], o_user_10_00_lut_03[15])
`ACX_BIND_USER_DESIGN_PORT(mcio_vio_oe[0], o_user_10_00_lut_03[8])
`ACX_BIND_USER_DESIGN_PORT(mcio_vio_oe[1], o_user_10_00_lut_03[9])
`ACX_BIND_USER_DESIGN_PORT(mcio_vio_oe[2], o_user_10_00_lut_03[10])
`ACX_BIND_USER_DESIGN_PORT(mcio_vio_oe[3], o_user_10_00_lut_03[11])
`ACX_BIND_USER_DESIGN_PORT(mcio_vio_out[0], o_user_10_00_lut_04[4])
`ACX_BIND_USER_DESIGN_PORT(mcio_vio_out[1], o_user_10_00_lut_04[12])
`ACX_BIND_USER_DESIGN_PORT(mcio_vio_out[2], o_user_10_00_lut_04[20])
`ACX_BIND_USER_DESIGN_PORT(mcio_vio_out[3], o_user_10_00_lut_05[0])
`ACX_BIND_USER_DESIGN_PORT(test[2], o_user_10_00_lut_03[24])
`ACX_BIND_USER_DESIGN_PORT(test_oe[2], o_user_10_00_lut_03[7])
`endif
    // Ports for vp_gpio_s_b2
`ifdef ACX_GPIO_S_FULL
    // Core Data
`ACX_BIND_USER_DESIGN_PORT(fpga_sys_scl_in, i_user_10_00_lut_01[21])
`ACX_BIND_USER_DESIGN_PORT(fpga_sys_sda_in, i_user_10_00_lut_02[1])
`ACX_BIND_USER_DESIGN_PORT(mcio_scl_in, i_user_10_00_lut_00[17])
`ACX_BIND_USER_DESIGN_PORT(mcio_sda_in, i_user_10_00_lut_00[25])
`ACX_BIND_USER_DESIGN_PORT(fpga_sys_scl_oe, o_user_10_00_lut_00[6])
`ACX_BIND_USER_DESIGN_PORT(fpga_sys_scl_out, o_user_10_00_lut_02[2])
`ACX_BIND_USER_DESIGN_PORT(fpga_sys_sda_oe, o_user_10_00_lut_00[7])
`ACX_BIND_USER_DESIGN_PORT(fpga_sys_sda_out, o_user_10_00_lut_02[10])
`ACX_BIND_USER_DESIGN_PORT(mcio_oe1_l, o_user_10_00_lut_01[14])
`ACX_BIND_USER_DESIGN_PORT(mcio_oe1_l_oe, o_user_10_00_lut_00[4])
`ACX_BIND_USER_DESIGN_PORT(mcio_oe_45_l, o_user_10_00_lut_01[22])
`ACX_BIND_USER_DESIGN_PORT(mcio_oe_45_l_oe, o_user_10_00_lut_00[5])
`ACX_BIND_USER_DESIGN_PORT(mcio_scl_oe, o_user_10_00_lut_00[2])
`ACX_BIND_USER_DESIGN_PORT(mcio_scl_out, o_user_10_00_lut_00[26])
`ACX_BIND_USER_DESIGN_PORT(mcio_sda_oe, o_user_10_00_lut_00[3])
`ACX_BIND_USER_DESIGN_PORT(mcio_sda_out, o_user_10_00_lut_01[6])
`endif
    // Ports for vp_pll_nw_2
`ifdef ACX_CLK_NW_FULL
`ACX_BIND_USER_DESIGN_PORT(pll_nw_2_ref0_312p5_clk, i_user_06_09_trunk_00[0])
`ACX_BIND_USER_DESIGN_PORT(vp_pll_nw_2_lock, i_user_00_08_lut_17[2])
`endif
    // Ports for vp_pll_sw_2
`ifdef ACX_CLK_SW_FULL
`ACX_BIND_USER_DESIGN_PORT(pll_sw_2_ref1_312p5_clk, i_user_06_00_trunk_00[3])
`ACX_BIND_USER_DESIGN_PORT(vp_pll_sw_2_lock, i_user_00_01_lut_17[2])
`endif

//////////////////////////////////////
// End IO Ring User Design Port Binding Include File
//////////////////////////////////////
