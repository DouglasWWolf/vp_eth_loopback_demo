//////////////////////////////////////
// ACE GENERATED VERILOG INCLUDE FILE
// Generated on: 2023.05.10 at 14:47:42 PDT
// By: ACE 9.0.1
// From project: vp_project
//////////////////////////////////////
// User Design Signal List Include File
//////////////////////////////////////

    // Ports for ethernet_0
    // Clocks and Resets
    logic        ethernet_0_m0_ff_clk_divby2;
    logic        ethernet_0_m1_ff_clk_divby2;
    logic        ethernet_0_ref_clk_divby2;
    // Free Running Counter
    logic  [63:0] ethernet_0_free_running_counter;
    // Quad MAC 0 Flow Control
    logic  [3:0] ethernet_0_quad0_emac_enable;
    logic  [3:0] ethernet_0_quad0_emac_pause_en;
    logic  [31:0] ethernet_0_quad0_emac_pause_on;
    logic  [31:0] ethernet_0_quad0_emac_xoff_gen;
    logic  [3:0] ethernet_0_quad0_lpi_txhold;
    logic  [3:0] ethernet_0_quad0_mac_stop_tx;
    logic  [3:0] ethernet_0_quad0_tx_hold_req;
    // Quad MAC 0 Status
    logic  [3:0] ethernet_0_m0_ffe_tx_ovr;
    logic  [3:0] ethernet_0_m0_ffp_tx_ovr;
    logic  [3:0] ethernet_0_m0_mac_tx_underflow;
    // Quad MAC 0 TSN
    logic  [255:0] ethernet_0_quad0_tx_ts;
    logic  [15:0] ethernet_0_quad0_tx_ts_id;
    logic  [3:0] ethernet_0_quad0_tx_ts_val;
    logic  [119:0] ethernet_0_quad0_peer_delay;
    logic  [3:0] ethernet_0_quad0_peer_delay_val;
    // Ports for noc
    // Ports for pll_ddr
    logic        pll_ddr_lock;
    // Ports for pll_eth_sys_ne_0
    logic        pll_eth_sys_ne_0_lock;
    // Ports for pll_gddr_SE
    logic        pll_gddr_SE_lock;
    // Ports for pll_gddr_SW
    logic        pll_gddr_SW_lock;
    // Ports for pll_noc_ne_1
    logic        i_clk;
    logic        i_eth_ts_clk;
    logic        i_reg_clk;
    logic        pll_noc_ne_1_lock;
    // Ports for pll_pcie
    logic        pll_pcie_lock;
    // Ports for vp_clkio_ne
    logic        fpga_rst_l;
    // Ports for vp_clkio_nw
    // Ports for vp_clkio_se
    // Ports for vp_clkio_sw
    // Ports for vp_gpio_n_b0
    // Core Data
    // Port name: ext_gpio_fpga_in[0] has been automatically combined into a the bussed signal below.
    logic        ext_gpio_fpga_in[7:0];
    // Port name: ext_gpio_fpga_in[1] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_in[2] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_in[3] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_in[4] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_in[5] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_in[6] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_in[7] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_oe[0] has been automatically combined into a the bussed signal below.
    logic        ext_gpio_fpga_oe[7:0];
    // Port name: ext_gpio_fpga_oe[1] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_oe[2] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_oe[3] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_oe[4] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_oe[5] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_oe[6] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_oe[7] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_out[0] has been automatically combined into a the bussed signal below.
    logic        ext_gpio_fpga_out[7:0];
    // Port name: ext_gpio_fpga_out[1] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_out[2] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_out[3] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_out[4] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_out[5] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_out[6] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_fpga_out[7] has been automatically combined into a bussed signal.
    logic        ext_gpio_oe_l;
    logic        ext_gpio_oe_l_oe;
    logic        led_oe_l;
    logic        led_oe_l_oe;
    // Ports for vp_gpio_n_b1
    // Core Data
    // Port name: ext_gpio_dir[0] has been automatically combined into a the bussed signal below.
    logic        ext_gpio_dir[7:0];
    // Port name: ext_gpio_dir[1] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir[2] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir[3] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir[4] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir[5] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir[6] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir[7] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir_oe[0] has been automatically combined into a the bussed signal below.
    logic        ext_gpio_dir_oe[7:0];
    // Port name: ext_gpio_dir_oe[1] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir_oe[2] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir_oe[3] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir_oe[4] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir_oe[5] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir_oe[6] has been automatically combined into a bussed signal.
    // Port name: ext_gpio_dir_oe[7] has been automatically combined into a bussed signal.
    // Port name: led_l[4] has been automatically combined into a the bussed signal below.
    logic        led_l[7:0];
    // Port name: led_l[5] has been automatically combined into a bussed signal.
    // Port name: led_l_oe[4] has been automatically combined into a the bussed signal below.
    logic        led_l_oe[7:0];
    // Port name: led_l_oe[5] has been automatically combined into a bussed signal.
    // Ports for vp_gpio_n_b2
    // Core Data
    // Port name: led_l[0] has been automatically combined into a bussed signal.
    // Port name: led_l[1] has been automatically combined into a bussed signal.
    // Port name: led_l[2] has been automatically combined into a bussed signal.
    // Port name: led_l[3] has been automatically combined into a bussed signal.
    // Port name: led_l[6] has been automatically combined into a bussed signal.
    // Port name: led_l[7] has been automatically combined into a bussed signal.
    // Port name: led_l_oe[0] has been automatically combined into a bussed signal.
    // Port name: led_l_oe[1] has been automatically combined into a bussed signal.
    // Port name: led_l_oe[2] has been automatically combined into a bussed signal.
    // Port name: led_l_oe[3] has been automatically combined into a bussed signal.
    // Port name: led_l_oe[6] has been automatically combined into a bussed signal.
    // Port name: led_l_oe[7] has been automatically combined into a bussed signal.
    // Ports for vp_gpio_s_b0
    // Core Data
    logic        fpga_avr_rxd;
    logic        fpga_ftdi_rxd;
    logic        fpga_i2c_mux_gnt;
    logic        irq_to_fpga;
    logic        qsfp_int_fpga_l;
    logic        fpga_avr_txd;
    logic        fpga_avr_txd_oe;
    logic        fpga_ftdi_txd;
    logic        fpga_ftdi_txd_oe;
    logic        fpga_i2c_req_l;
    logic        fpga_i2c_req_l_oe;
    logic        irq_to_avr;
    logic        irq_to_avr_oe;
    // Port name: test[1] has been automatically combined into a the bussed signal below.
    logic        test[2:1];
    // Port name: test_oe[1] has been automatically combined into a the bussed signal below.
    logic        test_oe[2:1];
    // Ports for vp_gpio_s_b1
    // Core Clock
    logic        mcio_vio_45_10_clk;
    // Core Data
    // Port name: mcio_vio_in[0] has been automatically combined into a the bussed signal below.
    logic        mcio_vio_in[3:0];
    // Port name: mcio_vio_in[1] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_in[2] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_in[3] has been automatically combined into a bussed signal.
    // Port name: mcio_dir[0] has been automatically combined into a the bussed signal below.
    logic        mcio_dir[3:0];
    // Port name: mcio_dir[1] has been automatically combined into a bussed signal.
    // Port name: mcio_dir[2] has been automatically combined into a bussed signal.
    // Port name: mcio_dir[3] has been automatically combined into a bussed signal.
    logic        mcio_dir_45;
    logic        mcio_dir_45_oe;
    // Port name: mcio_dir_oe[0] has been automatically combined into a the bussed signal below.
    logic        mcio_dir_oe[3:0];
    // Port name: mcio_dir_oe[1] has been automatically combined into a bussed signal.
    // Port name: mcio_dir_oe[2] has been automatically combined into a bussed signal.
    // Port name: mcio_dir_oe[3] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_oe[0] has been automatically combined into a the bussed signal below.
    logic        mcio_vio_oe[3:0];
    // Port name: mcio_vio_oe[1] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_oe[2] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_oe[3] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_out[0] has been automatically combined into a the bussed signal below.
    logic        mcio_vio_out[3:0];
    // Port name: mcio_vio_out[1] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_out[2] has been automatically combined into a bussed signal.
    // Port name: mcio_vio_out[3] has been automatically combined into a bussed signal.
    // Port name: test[2] has been automatically combined into a bussed signal.
    // Port name: test_oe[2] has been automatically combined into a bussed signal.
    // Ports for vp_gpio_s_b2
    // Core Data
    logic        fpga_sys_scl_in;
    logic        fpga_sys_sda_in;
    logic        mcio_scl_in;
    logic        mcio_sda_in;
    logic        fpga_sys_scl_oe;
    logic        fpga_sys_scl_out;
    logic        fpga_sys_sda_oe;
    logic        fpga_sys_sda_out;
    logic        mcio_oe1_l;
    logic        mcio_oe1_l_oe;
    logic        mcio_oe_45_l;
    logic        mcio_oe_45_l_oe;
    logic        mcio_scl_oe;
    logic        mcio_scl_out;
    logic        mcio_sda_oe;
    logic        mcio_sda_out;
    // Ports for vp_pll_nw_2
    logic        pll_nw_2_ref0_312p5_clk;
    logic        vp_pll_nw_2_lock;
    // Ports for vp_pll_sw_2
    logic        pll_sw_2_ref1_312p5_clk;
    logic        vp_pll_sw_2_lock;

//////////////////////////////////////
// End User Design Signal List Include File
//////////////////////////////////////
